library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package spi_master_pkg is
  constant spi_num_bits : positive := 8; 
end package;

package body spi_master_pkg is
end package body;